//-------------------------------------------------------------------------------------------------
module rom
//-------------------------------------------------------------------------------------------------
#
(
        parameter KB = 0
)
(
        input  wire                      clock,
        input  wire[$clog2(KB*1024)-1:0] address,
        output reg [                7:0] q
);
//-------------------------------------------------------------------------------------------------

reg[7:0] rom[(KB*1024)-1:0];
always @(posedge clock)  q <= rom[a];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------